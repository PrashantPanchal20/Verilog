module and_gate_data_flow(a,b,c);
    input a;
    input b;
    output c;

assign c = a & b ;

endmodule
